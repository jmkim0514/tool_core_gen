module slave (
    input             i_clk,
    input             i_valid,
    output            o_ready

);

endmodule