module crm (
    input                   i_xin   ,
    input                   i_por   ,
    output                  o_clk_100,
    output                  o_clk_200,
    output                  o_clk_300,
    output                  o_clk_600,
    output                  o_clk_100,
    output                  o_clk_200,
    output                  o_clk_300,
    output                  o_clk_600,
    output                  o_rstn_100,
    output                  o_rstn_200,
    output                  o_rstn_300,
    output                  o_rstn_600,
    output                  o_rstn_100,
    output                  o_rstn_200,
    output                  o_rstn_300,
    output                  o_rstn_600
);


endmodule