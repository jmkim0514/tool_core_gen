module crm (
    input             i_clk,
    output            o_clk_mst,
    output            o_clk_slv

);

endmodule