module crm_peri (
    input           i_clk_100,
    input           i_rstn_100,
    
    output          o_clk_ssp,
    output          o_rstn_ssp,
    output          o_clk_gpio,
    output          o_rstn_gpio,
    output          o_clk_i2c,
    output          o_rstn_i2c

);


endmodule