module master (
    input             i_clk,
    output            o_mst_valid,
    input             i_mst_ready

);

endmodule