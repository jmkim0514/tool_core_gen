module crm (
    input                   i_xin   ,
    output                  o_pclk   ,
    output                  o_hclk   ,
    output                  o_xclk   ,
    output                  o_presetn,
    output                  o_hresetn,
    output                  o_xresetn,
    output                  o_irq    ,
    input                   i_irq
);


endmodule