module crm_cpu (
    input           i_clk_200,
    input           i_clk_100,
    input           i_rstn_200,
    input           i_rstn_100,
    
    output          o_clk_cpu,
    output          o_clk_peri,
    output          o_rstn_cpu,
    output          o_rstn_peri
);


endmodule